-- fpga_config.vhd: user constants
use work.clkgen_cfg.all;

package fpga_cfg is
   constant DCM_FREQUENCY : dcm_freq := DCM_40MHz;
end fpga_cfg;

package body fpga_cfg is
end fpga_cfg;
